library verilog;
use verilog.vl_types.all;
entity tb_led is
end tb_led;
